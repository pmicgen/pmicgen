.subckt ota
M5 id  id vss vss sky130_fd_pr__nfet_01v8 L= W= nf= stack=
.ends ota